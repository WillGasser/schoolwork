library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity test_decoder is
end test_decoder;

architecture Behavioral of test_decoder is
  component twobitdecoder is
    generic(prop_delay: time := 10 ns);
    port(
      encoded: in bit_vector(1 downto 0);
      out0, out1, out2, out3: out bit
    );
  end component;
  signal encoded: bit_vector(1 downto 0) := "00";
  signal out0, out1, out2, out3: bit;
begin
  uut: twobitdecoder
    generic map(prop_delay => 10 ns)
    port map(
      encoded => encoded,
      out0 => out0,
      out1 => out1,
      out2 => out2,
      out3 => out3
    );
  process
  begin
    encoded <= "00"; wait for 20 ns;
    encoded <= "01"; wait for 20 ns;
    encoded <= "10"; wait for 20 ns;
    encoded <= "11"; wait for 20 ns;
    wait;
  end process;
end Behavioral;
